-------------------------------------------------------------------------------
-- Engineer:       Berger Jonas
-- Create Date:    2024-10-05
-- Design Name:    Dummy Value Generater
-- Module Name:    dummy_gen - rtl
-- Project Name:   Sensor Actuator Emulator
-- Revision:       v1.0
-------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity imu_sensor_dummy_gen is
  generic (
    G_IMU_DATA_CNT : natural := 500
  );
  port (
    clk_i  : in std_logic;
    rst_i  : in std_logic;
    tick_i : in std_logic;

    accel_xout_o : out std_logic_vector(15 downto 0);
    accel_yout_o : out std_logic_vector(15 downto 0);
    accel_zout_o : out std_logic_vector(15 downto 0);
    gyro_xout_o  : out std_logic_vector(15 downto 0);
    gyro_yout_o  : out std_logic_vector(15 downto 0);
    gyro_zout_o  : out std_logic_vector(15 downto 0);
    mag_xout_o   : out std_logic_vector(15 downto 0);
    mag_yout_o   : out std_logic_vector(15 downto 0);
    mag_zout_o   : out std_logic_vector(15 downto 0);
    temp_out_o   : out std_logic_vector(15 downto 0)
  );
end entity imu_sensor_dummy_gen;

architecture rtl of imu_sensor_dummy_gen is

  type dummy_lut_t is array (0 to G_IMU_DATA_CNT-1) of std_logic_vector(15 downto 0);

  signal s_dummy_accelx_lut : dummy_lut_t := (
  x"FFD2", x"FFD9", x"FFD6", x"FFD9", x"FF67", x"0031", x"FFD2", x"FFE0",
  x"FFAA", x"FF7E", x"0011", x"FFA1", x"FF51", x"FFB9", x"FFED", x"FFBF",
  x"FF68", x"0FFF", x"FF31", x"FF6E", x"FF5B", x"FF5E", x"FFBF", x"FFDE",
  x"FFE4", x"FF2F", x"0034", x"FFCB", x"000F", x"0012", x"0026", x"001D",
  x"002F", x"003A", x"0037", x"0095", x"006E", x"0081", x"00A7", x"00DC",
  x"015D", x"011A", x"00CA", x"0173", x"01C3", x"01D0", x"01F5", x"002F",
  x"0226", x"0213", x"028C", x"02D4", x"02E0", x"003E", x"02F9", x"0315",
  x"032F", x"037F", x"03BE", x"03C8", x"039F", x"03E6", x"03DB", x"03CF",
  x"03F2", x"03FB", x"0410", x"0040", x"0433", x"0435", x"041D", x"0423",
  x"042D", x"0430", x"0452", x"044B", x"0442", x"0428", x"042E", x"0046",
  x"03A5", x"03BD", x"03A0", x"03AE", x"038B", x"03BC", x"03EB", x"03AF",
  x"0387", x"03B8", x"03BA", x"03C6", x"019D", x"02BE", x"032F", x"0342",
  x"02FC", x"0297", x"022E", x"0192", x"0183", x"018B", x"013A", x"00DF",
  x"00BC", x"0095", x"0071", x"00B9", x"00D6", x"00B2", x"00BB", x"0099",
  x"00A5", x"00EB", x"001B", x"00BB", x"00A8", x"00B6", x"00D7", x"00B2",
  x"0091", x"0084", x"0087", x"008D", x"0061", x"006A", x"0061", x"FFBC",
  x"FF9A", x"FFA3", x"FFB8", x"FFCE", x"FFC2", x"003F", x"FFE3", x"FF8D",
  x"FF67", x"FF4D", x"FF5B", x"FF9C", x"FEA2", x"FECA", x"FD69", x"FD47",
  x"FD67", x"FE1D", x"FE17", x"0FE7", x"FE6D", x"0FF6", x"FFBE", x"0064",
  x"00B4", x"00CE", x"0115", x"014C", x"019E", x"01CD", x"01D5", x"019E",
  x"01BE", x"01E6", x"01CA", x"01A3", x"01AD", x"0164", x"01C7", x"01ED",
  x"01D0", x"0184", x"014F", x"0011", x"00AE", x"0039", x"FF56", x"FF7B",
  x"FFC5", x"FFEB", x"FF82", x"FEA1", x"FEAB", x"FE99", x"FE80", x"0FE0",
  x"FD55", x"FCCE", x"0FD0", x"FCFD", x"FCF6", x"FCAF", x"0FCF", x"FBAA",
  x"FBCE", x"FBC6", x"FB89", x"FB8D", x"FAFF", x"FA68", x"FA45", x"FA24",
  x"FA19", x"F9B6", x"F959", x"F923", x"F92A", x"F932", x"0F9E", x"F91C",
  x"F92A", x"F944", x"F947", x"F8FE", x"F8A6", x"F826", x"F7F3", x"F841",
  x"F84C", x"F830", x"F85D", x"F899", x"F8B8", x"F885", x"F949", x"F9BF",
  x"F9FF", x"F98E", x"F9A7", x"0FA0", x"FA2B", x"FA6B", x"FAD5", x"FB17",
  x"FB6B", x"FBC6", x"FC3C", x"FCB8", x"FD5C", x"FDF5", x"FE65", x"FE90",
  x"FE89", x"FED4", x"FEBE", x"FF58", x"FFE1", x"0019", x"0032", x"005A",
  x"009C", x"00C5", x"014E", x"0189", x"01B2", x"0226", x"0243", x"002C",
  x"021F", x"0272", x"02CE", x"003E", x"0341", x"0343", x"0379", x"03B4",
  x"03FC", x"043F", x"043D", x"004F", x"03DC", x"03F8", x"043A", x"041A",
  x"004B", x"0434", x"0488", x"04DE", x"005F", x"0531", x"057F", x"05A5",
  x"0589", x"059A", x"05A4", x"0580", x"0566", x"0554", x"053E", x"054E",
  x"056E", x"0056", x"04AE", x"0456", x"0412", x"004D", x"03D1", x"0364",
  x"0339", x"02EF", x"0291", x"0253", x"024E", x"0249", x"0224", x"002F",
  x"01A5", x"01A2", x"0188", x"015A", x"017F", x"0142", x"00C2", x"000D",
  x"FFF9", x"002B", x"0025", x"FFED", x"FF96", x"FF56", x"FF34", x"FF59",
  x"FF93", x"FF6D", x"FF33", x"FF32", x"FF3B", x"FF3C", x"FF53", x"FF4F",
  x"FF79", x"FFA3", x"FF86", x"FF93", x"FF9C", x"FFC7", x"FFFB", x"FFE0",
  x"0018", x"003B", x"003F", x"0049", x"0066", x"0038", x"0030", x"0021",
  x"FFFD", x"FFE9", x"FFF5", x"003D", x"001C", x"FFF1", x"FFCE", x"FFB2",
  x"FFD2", x"FFD3", x"FFF2", x"FFE6", x"FFB1", x"FFA5", x"FF9D", x"FF60",
  x"FF3A", x"FF4D", x"FF8B", x"FFA9", x"FF77", x"FF69", x"FF63", x"FF93",
  x"FF54", x"FF47", x"FF5B", x"FF3A", x"FF17", x"FF17", x"0FF7", x"FF14",
  x"FF1D", x"FF13", x"0FF7", x"FEF4", x"FEE4", x"FF49", x"FF77", x"FFC2",
  x"FFAD", x"FFA0", x"FFAF", x"FFB6", x"FFE4", x"002C", x"001F", x"FFE4",
  x"FFD0", x"004A", x"0020", x"006C", x"006C", x"004F", x"007F", x"00AD",
  x"00EF", x"00EC", x"00B2", x"00AF", x"005C", x"001A", x"005E", x"009E",
  x"00B3", x"0050", x"003F", x"FFDD", x"0087", x"0038", x"0069", x"0038",
  x"FFFB", x"FFF9", x"002E", x"005A", x"0026", x"002C", x"0004", x"FFD7",
  x"FFFF", x"FFC4", x"FFDD", x"FFE5", x"0015", x"000D", x"0000", x"FFF8",
  x"FFFA", x"0000", x"0048", x"0077", x"00A5", x"0081", x"0050", x"00C7",
  x"00A5", x"00AC", x"00C6", x"0015", x"0015", x"00DB", x"00DA", x"00CE",
  x"00BD", x"00CA", x"00C0", x"0087", x"009C", x"00FC", x"0112", x"00F0",
  x"00A9", x"0076", x"0075", x"0069", x"0094", x"007E", x"0036", x"001F",
  x"000F", x"FFFA", x"0017", x"0025", x"0036", x"0058", x"0021", x"0049",
  x"0097", x"00E4", x"00FE", x"00B5", x"00C6", x"00E9", x"001E", x"0133",
  x"019B", x"01E0", x"01C0", x"01C7", x"01F6", x"0221", x"0271", x"02D3",
  x"02C3", x"02DC", x"0343", x"035C", x"0366", x"03CD", x"0432", x"0495",
  x"0496", x"04A0", x"0056", x"052E"
  );

  signal s_dummy_accely_lut : dummy_lut_t := (
  x"FFC5", x"FFBE", x"FFB0", x"FFB8", x"FF9C", x"FFCB", x"FFB9", x"FFA4",
  x"FFB9", x"FFAB", x"FFD3", x"FFCF", x"FFFA", x"FF97", x"FFE1", x"001E",
  x"0042", x"FF4F", x"FFB8", x"FF6B", x"FFDA", x"003D", x"0071", x"00DE",
  x"0017", x"FDEF", x"016E", x"0072", x"00FE", x"0151", x"012F", x"019B",
  x"0253", x"02C9", x"028B", x"028C", x"029E", x"0363", x"004B", x"03E1",
  x"0442", x"04B8", x"04B2", x"03EA", x"046D", x"04C3", x"0436", x"0530",
  x"05D3", x"0041", x"03E0", x"0444", x"0041", x"03B8", x"038E", x"02D8",
  x"01ED", x"001F", x"00F0", x"0119", x"00B3", x"0093", x"00B8", x"007A",
  x"0078", x"0018", x"FF5C", x"FEA2", x"FEE6", x"0FF7", x"FFD8", x"FFC1",
  x"FE61", x"FD92", x"FDCD", x"FEE1", x"0FF4", x"FF52", x"0FF1", x"FE24",
  x"FD1B", x"FB8B", x"FB51", x"FBFB", x"FC50", x"FC61", x"FCA3", x"FC9E",
  x"FC34", x"FC5D", x"FC48", x"FC50", x"FC38", x"FB21", x"FB47", x"FB4C",
  x"FB8A", x"FBF1", x"FC60", x"FC86", x"FC3D", x"FC74", x"FD18", x"FD7A",
  x"FD83", x"FD8C", x"FD7B", x"FD94", x"FE32", x"FE25", x"FE3F", x"FE4B",
  x"FE32", x"FE52", x"FE14", x"FE60", x"FEC4", x"FE93", x"FED6", x"0FFC",
  x"FEFC", x"FF50", x"FF55", x"FF6A", x"FF53", x"FFB4", x"FED8", x"FE44",
  x"FF4D", x"FF65", x"FFD8", x"FFDA", x"0055", x"FF98", x"FFFE", x"000B",
  x"005F", x"0009", x"FFEF", x"FF98", x"FF11", x"0FFA", x"FD1E", x"FC9E",
  x"FDCA", x"FEC6", x"FF81", x"004E", x"00C4", x"011F", x"0144", x"01DC",
  x"0276", x"02B4", x"02A5", x"02F6", x"02DB", x"003A", x"02F6", x"02CC",
  x"0031", x"02C3", x"0295", x"029B", x"0261", x"01D9", x"01B5", x"0166",
  x"00B6", x"0044", x"0030", x"0097", x"00A3", x"0086", x"008E", x"0053",
  x"004F", x"FFFC", x"FF76", x"FFB1", x"FFCF", x"FFC4", x"FFA8", x"FF81",
  x"FFB6", x"0040", x"0076", x"006B", x"FFCB", x"FF83", x"FF40", x"FF77",
  x"FFB1", x"FFE0", x"0008", x"000D", x"0042", x"FFEC", x"FF96", x"FFC5",
  x"FFF3", x"FFA3", x"FFB3", x"FFC3", x"FFD3", x"FFCC", x"FFF7", x"000F",
  x"FFE8", x"FFB5", x"FF74", x"FF6E", x"FFC2", x"FFEC", x"FFF6", x"0057",
  x"0022", x"FFD7", x"FF89", x"FF83", x"FFA2", x"FF6E", x"FFF6", x"004C",
  x"0066", x"00D3", x"00BE", x"004E", x"FFE6", x"FF1E", x"FFBC", x"FFDA",
  x"FFFA", x"002F", x"0053", x"00C4", x"00AC", x"001B", x"0023", x"004E",
  x"0055", x"0009", x"0019", x"0023", x"0092", x"001A", x"00F0", x"0099",
  x"00D0", x"0146", x"0188", x"0169", x"0136", x"0138", x"0012", x"0122",
  x"0143", x"012C", x"00FA", x"00E5", x"012F", x"0180", x"01A8", x"01A6",
  x"0191", x"01C2", x"01BE", x"01AE", x"01FD", x"01FF", x"01FF", x"01B2",
  x"01C6", x"01D0", x"01DC", x"0029", x"002B", x"025B", x"028A", x"02A3",
  x"027A", x"0219", x"021C", x"0234", x"0231", x"0235", x"01F4", x"01ED",
  x"01F6", x"01E1", x"0020", x"0244", x"0252", x"023A", x"019F", x"0115",
  x"00DC", x"0098", x"00A1", x"00EC", x"00A0", x"005B", x"0085", x"00B4",
  x"00D7", x"00D3", x"00BE", x"0053", x"002C", x"0084", x"002F", x"FFE7",
  x"FFD6", x"FF8B", x"FF96", x"FF9F", x"FF6E", x"FF5E", x"FF37", x"FF1E",
  x"FF1F", x"FF11", x"FECD", x"FEC5", x"FEF5", x"FF60", x"FF68", x"FF40",
  x"FF2F", x"FF40", x"FF2D", x"FF23", x"0FF9", x"FEBB", x"FE5A", x"FE59",
  x"FE3C", x"FE23", x"FDD6", x"FD87", x"FD45", x"FCEE", x"FCB4", x"FC80",
  x"FC27", x"FBBE", x"FBC6", x"FBDC", x"FBCE", x"FAF4", x"0FB2", x"FACC",
  x"FA9F", x"FA67", x"FA88", x"FA51", x"F9C9", x"F98A", x"F95B", x"F8D5",
  x"F894", x"F87E", x"F8AF", x"F899", x"F87B", x"F826", x"0F8B", x"F83D",
  x"F7B3", x"F7A7", x"F7BE", x"F7B3", x"F76D", x"F751", x"F763", x"F775",
  x"F784", x"F74B", x"F769", x"F7A7", x"F7E1", x"F7D7", x"F858", x"F921",
  x"F96B", x"F95E", x"F977", x"F99D", x"F9AC", x"F9F3", x"FA57", x"FAE7",
  x"FB42", x"FBD2", x"FBBC", x"FC6C", x"FD26", x"FD7B", x"FDA4", x"FE4E",
  x"0FF6", x"FFBA", x"FF8E", x"FF84", x"FF54", x"FFA1", x"0091", x"0119",
  x"0125", x"00EB", x"00FA", x"014B", x"0195", x"0310", x"035E", x"0379",
  x"0332", x"0359", x"03F0", x"04BA", x"04D8", x"04D8", x"0522", x"0570",
  x"0583", x"0583", x"0562", x"0583", x"062A", x"0658", x"0061", x"05FF",
  x"061A", x"066B", x"067B", x"06A2", x"06FA", x"0731", x"075D", x"07BE",
  x"07DC", x"0822", x"008F", x"07C8", x"0830", x"085E", x"0853", x"0852",
  x"0856", x"089B", x"086F", x"0824", x"07C1", x"0765", x"072A", x"0721",
  x"06AB", x"061D", x"05E1", x"05D1", x"05F9", x"05DA", x"0577", x"005E",
  x"04D9", x"0460", x"03EB", x"035F", x"02C9", x"0266", x"0227", x"01D4",
  x"0015", x"0087", x"0049", x"009D", x"00B1", x"00CB", x"00B8", x"00A1",
  x"0090", x"0073", x"009A", x"004B", x"FFFE", x"0000", x"0060", x"00EB",
  x"00EE", x"0094", x"00F6", x"0114", x"00F3", x"001F", x"0142", x"0260",
  x"0024", x"0149", x"0135", x"0184"
  );

  signal s_dummy_accelz_lut : dummy_lut_t := (
  x"0086", x"07FA", x"07FD", x"07F2", x"0081", x"008D", x"0087", x"008D",
  x"008D", x"0083", x"07FF", x"008F", x"008A", x"0819", x"0864", x"0840",
  x"081D", x"08EC", x"0A34", x"098A", x"0828", x"077A", x"07C2", x"07C6",
  x"08F8", x"08E2", x"084D", x"07C3", x"07A5", x"07D0", x"0819", x"07D2",
  x"07A0", x"07F3", x"07FF", x"07FA", x"078F", x"06EA", x"06A7", x"06CB",
  x"0699", x"06E4", x"06D7", x"056F", x"05D8", x"0670", x"05A7", x"0593",
  x"0694", x"063A", x"0525", x"0537", x"0622", x"06FE", x"06BE", x"05FC",
  x"0523", x"0585", x"06BC", x"0780", x"075A", x"06EA", x"06BD", x"0676",
  x"0632", x"0660", x"0073", x"079B", x"06B1", x"06A3", x"05FD", x"0069",
  x"05FB", x"064A", x"0698", x"062E", x"05BF", x"05D2", x"0584", x"0636",
  x"06D0", x"079D", x"0747", x"0681", x"069E", x"0671", x"05B2", x"0610",
  x"0554", x"05A3", x"0617", x"06A7", x"0678", x"0692", x"066F", x"073D",
  x"074B", x"0749", x"0723", x"0728", x"06F9", x"06FD", x"07AD", x"07DA",
  x"07DC", x"0087", x"082D", x"008F", x"0081", x"0086", x"0774", x"072B",
  x"076F", x"0770", x"071E", x"06ED", x"071A", x"0753", x"07B0", x"07A0",
  x"0784", x"07D8", x"07D7", x"0845", x"0854", x"0082", x"08B3", x"0836",
  x"081A", x"07FA", x"07B8", x"0818", x"07E3", x"0823", x"0789", x"0818",
  x"0895", x"0089", x"07E8", x"07D9", x"085B", x"0798", x"0A3E", x"0A7F",
  x"07D3", x"0769", x"087D", x"091D", x"094D", x"08C2", x"07BF", x"06CA",
  x"0076", x"077F", x"0757", x"06D4", x"06D1", x"0077", x"072E", x"078F",
  x"07F9", x"0816", x"07F9", x"07AD", x"0739", x"07BA", x"0676", x"06B9",
  x"0694", x"06FA", x"06FD", x"072F", x"0725", x"076E", x"0854", x"0868",
  x"078F", x"06F0", x"007B", x"07B8", x"078C", x"078C", x"0747", x"06B9",
  x"07CC", x"081B", x"07D4", x"073A", x"06B5", x"0632", x"06A3", x"0077",
  x"065D", x"0068", x"0638", x"05BA", x"05A4", x"0614", x"061A", x"05D4",
  x"0570", x"0576", x"05D1", x"05B9", x"0528", x"053A", x"0563", x"005F",
  x"04A5", x"047B", x"043C", x"0477", x"04DB", x"0589", x"05C0", x"051D",
  x"0056", x"0565", x"0561", x"0563", x"0577", x"059C", x"055B", x"04EF",
  x"0567", x"0657", x"06C4", x"06B4", x"06AD", x"061E", x"0656", x"06AA",
  x"0072", x"0718", x"06F8", x"06B3", x"0657", x"06B2", x"0075", x"0742",
  x"077C", x"0785", x"0753", x"074D", x"0743", x"0721", x"0746", x"07B6",
  x"0872", x"0837", x"077A", x"073E", x"0757", x"0736", x"072E", x"07D7",
  x"0814", x"07AA", x"071B", x"06F4", x"06E0", x"072D", x"06FE", x"06B6",
  x"0658", x"05DB", x"05F4", x"0655", x"0714", x"06DE", x"0669", x"069A",
  x"06F0", x"068C", x"006D", x"0580", x"0540", x"0538", x"04E1", x"04A4",
  x"04F3", x"04C2", x"04AB", x"0511", x"0543", x"055E", x"059E", x"051D",
  x"0050", x"0551", x"05AD", x"064F", x"06C6", x"06B3", x"0681", x"06CF",
  x"069F", x"06A6", x"0758", x"07D5", x"078C", x"0077", x"074E", x"0761",
  x"07C1", x"07C3", x"07B8", x"07B6", x"0727", x"0713", x"07B0", x"08A9",
  x"08D0", x"07D4", x"0782", x"008A", x"0881", x"0893", x"08C8", x"0873",
  x"07E3", x"07F7", x"0852", x"0880", x"0881", x"0893", x"08B3", x"088E",
  x"0861", x"0833", x"0844", x"0850", x"0852", x"0088", x"0080", x"07C4",
  x"07B4", x"074E", x"0728", x"074E", x"0718", x"06E3", x"007B", x"0721",
  x"06EF", x"0714", x"06E9", x"0654", x"0635", x"0667", x"068C", x"0653",
  x"05FC", x"05B4", x"054D", x"04F7", x"04FB", x"04F4", x"042F", x"042A",
  x"0047", x"03D9", x"034F", x"0031", x"02E8", x"0311", x"02C4", x"026A",
  x"0237", x"0229", x"0022", x"01E4", x"01FA", x"0023", x"01FD", x"0218",
  x"0020", x"023E", x"0284", x"02D1", x"0324", x"039B", x"0334", x"038A",
  x"0427", x"04B1", x"04FB", x"04F6", x"0535", x"04E9", x"04B3", x"0550",
  x"0626", x"06DA", x"06DA", x"0659", x"05F9", x"06DA", x"07D4", x"07CB",
  x"0759", x"06F2", x"0774", x"0795", x"07B2", x"008E", x"0081", x"079F",
  x"076F", x"075C", x"077D", x"07BC", x"0087", x"0719", x"0714", x"06F0",
  x"074B", x"0748", x"06CA", x"063E", x"006E", x"065F", x"0653", x"0626",
  x"0626", x"062A", x"05E5", x"053B", x"051B", x"053A", x"0541", x"04E5",
  x"04A7", x"0461", x"0049", x"03BC", x"039E", x"0363", x"0337", x"0284",
  x"025F", x"029E", x"0282", x"0028", x"01F0", x"024E", x"026D", x"0282",
  x"029A", x"02C9", x"02D7", x"0315", x"0333", x"0353", x"0348", x"0370",
  x"03D7", x"0448", x"04C9", x"04FD", x"051A", x"053B", x"059F", x"0633",
  x"06DF", x"0744", x"074D", x"0749", x"06F4", x"073A", x"07FB", x"085D",
  x"07A8", x"06D0", x"06A0", x"07F3", x"08F1", x"08D0", x"084F", x"008E",
  x"07DF", x"07BA", x"0811", x"0832", x"07C6", x"0754", x"0747", x"0733",
  x"071B", x"072F", x"06CF", x"068F", x"072D", x"0681", x"05F1", x"06D0",
  x"0689", x"065F", x"0544", x"04DC"
  );

  signal s_dummy_gyrox_lut : dummy_lut_t := (
  x"FFF5", x"FFF5", x"FFEE", x"FFF7", x"FFDD", x"0020", x"0019", x"0007",
  x"0001", x"002F", x"0042", x"0041", x"0079", x"0084", x"009A", x"0032",
  x"000C", x"0057", x"00E3", x"01CF", x"02DC", x"0285", x"02A7", x"03A4",
  x"03E6", x"03FD", x"04BE", x"02CC", x"032A", x"0372", x"03B9", x"0491",
  x"0610", x"068A", x"008A", x"094E", x"093F", x"07EF", x"073A", x"05EA",
  x"0462", x"0392", x"03A8", x"0330", x"027A", x"00D5", x"FFC8", x"FF35",
  x"FE88", x"FE2E", x"FD66", x"FB9E", x"F961", x"F8B9", x"F88F", x"F886",
  x"F859", x"F841", x"F792", x"F844", x"F975", x"FB2D", x"FB75", x"FAD6",
  x"FA43", x"0FAD", x"FB2E", x"FC16", x"FDD2", x"FDEB", x"FDC9", x"FD65",
  x"FE57", x"FF6F", x"0011", x"0038", x"FFD7", x"FF47", x"FEFE", x"FE28",
  x"FDAE", x"FD9F", x"FF2E", x"FEF7", x"FEEF", x"FF93", x"FF98", x"FEF4",
  x"FE2C", x"0FE6", x"FD44", x"0FC5", x"FCA3", x"FDA8", x"00E1", x"0018",
  x"02C0", x"0434", x"03CA", x"03B4", x"03D1", x"0470", x"004A", x"03F3",
  x"0368", x"0358", x"035E", x"03CC", x"034D", x"0291", x"025B", x"01DD",
  x"01C2", x"025B", x"02EC", x"036E", x"02F7", x"0368", x"039E", x"038E",
  x"035A", x"0315", x"02E5", x"025B", x"0281", x"007C", x"0FFF", x"0063",
  x"02D6", x"031F", x"01EB", x"01A3", x"0087", x"00D1", x"0085", x"00EB",
  x"00B7", x"0112", x"00BB", x"00CC", x"008E", x"0143", x"00F7", x"000E",
  x"01B6", x"02FC", x"0324", x"031C", x"02E8", x"026C", x"0215", x"02A1",
  x"0248", x"0167", x"00C8", x"00E2", x"003B", x"000E", x"0005", x"FFE0",
  x"FF55", x"FE1E", x"FCEC", x"FC54", x"FBDD", x"FBEE", x"FC58", x"FCFC",
  x"0FD5", x"FCDF", x"FCC1", x"FCCA", x"FD1E", x"FDA5", x"FE12", x"FE3B",
  x"0FF0", x"FFC5", x"FFE3", x"0034", x"000B", x"002E", x"0048", x"FFCE",
  x"FFF8", x"000C", x"0030", x"0029", x"0001", x"0059", x"00A1", x"0006",
  x"FFC5", x"FFE5", x"FFB3", x"0013", x"0058", x"0035", x"FFF4", x"FFF1",
  x"0019", x"FFD5", x"FFC3", x"FFD2", x"000E", x"FFA9", x"FF6D", x"FFCE",
  x"0006", x"002D", x"0051", x"FFE0", x"FFBB", x"FFAF", x"0024", x"005F",
  x"0048", x"003D", x"0085", x"00DD", x"00A4", x"007B", x"0064", x"003A",
  x"FF4D", x"FF4C", x"00E7", x"019D", x"01E5", x"00E9", x"005C", x"FFFC",
  x"004C", x"0076", x"00D8", x"01BD", x"025A", x"0188", x"0006", x"FF46",
  x"FF21", x"FFAF", x"000E", x"003A", x"FFED", x"0123", x"01FA", x"0185",
  x"00DF", x"0116", x"001E", x"01AE", x"002D", x"01BE", x"0156", x"0117",
  x"01B3", x"02AF", x"025F", x"0015", x"00F1", x"01B8", x"024D", x"0025",
  x"0120", x"00FA", x"00B1", x"00CD", x"015D", x"0175", x"00F0", x"00E6",
  x"0176", x"0233", x"0283", x"0218", x"01D1", x"01A5", x"0128", x"00B4",
  x"FFC6", x"FEC1", x"FE7C", x"FEB0", x"FEE8", x"FEEC", x"FE9D", x"FE78",
  x"FE2B", x"FDDC", x"FD57", x"FC3A", x"FB66", x"FB6C", x"FBC8", x"FBDD",
  x"0FC4", x"FC56", x"FC19", x"FC62", x"FD2E", x"FDE8", x"FDA0", x"FD64",
  x"FCF9", x"FD80", x"FDF4", x"FE78", x"FE77", x"FE5E", x"FE28", x"FD8B",
  x"FD1F", x"FD7A", x"FDB4", x"FD4B", x"FD3B", x"FD8A", x"FE1C", x"FEB6",
  x"FF37", x"FFA1", x"FFA4", x"FF68", x"FF7B", x"FFAF", x"FF7B", x"0FF8",
  x"FE37", x"FD3F", x"FCBD", x"FC64", x"FBFF", x"FB89", x"FA7B", x"FA57",
  x"FA28", x"F9DB", x"FB27", x"FB12", x"FA33", x"0FAF", x"F9F1", x"FA36",
  x"FAB7", x"FA7A", x"FA1F", x"FA1F", x"FA2B", x"F9DF", x"F9C5", x"F9C4",
  x"F988", x"F929", x"F955", x"F91E", x"F8B3", x"F8E0", x"F981", x"F9AE",
  x"F95F", x"F8D4", x"F98B", x"F9DD", x"FA72", x"FB42", x"FBBF", x"FCEB",
  x"FD53", x"FD5C", x"FE20", x"FF4D", x"0016", x"00C2", x"0221", x"0037",
  x"0355", x"03AF", x"0556", x"066E", x"0748", x"07B6", x"079D", x"0726",
  x"075E", x"0798", x"07AD", x"088E", x"08A6", x"083C", x"07EE", x"0973",
  x"0C78", x"0B6F", x"0ADF", x"09E8", x"0A6C", x"0B26", x"0A3D", x"092E",
  x"0828", x"0829", x"0854", x"0840", x"0877", x"0846", x"0822", x"07BC",
  x"0752", x"0746", x"0785", x"0813", x"07B2", x"008B", x"0863", x"0856",
  x"07F2", x"07CD", x"075C", x"0756", x"06C1", x"0065", x"05D1", x"05D4",
  x"05BB", x"05E2", x"05B9", x"05C3", x"05A3", x"05F3", x"0064", x"0635",
  x"0683", x"06FB", x"0720", x"0768", x"0720", x"0635", x"05C2", x"04C7",
  x"03A6", x"02E3", x"0263", x"01DA", x"00DE", x"002E", x"FF64", x"FEDC",
  x"FD9E", x"FC44", x"FAE1", x"F9DA", x"F92E", x"F89A", x"F7E8", x"F768",
  x"0F71", x"F662", x"F5D5", x"F59C", x"F545", x"F4ED", x"F4BE", x"F4C7",
  x"F517", x"F54F", x"F569", x"F624", x"F780", x"F828", x"F8AE", x"FA86",
  x"FCB6", x"FDEA", x"FCA8", x"FB9A", x"FC3A", x"FD76", x"FEBF", x"FF4F",
  x"000B", x"FFBD", x"FF82", x"00D9", x"001C", x"016D", x"0176", x"0015",
  x"0043", x"0078", x"0133", x"00C3", x"00BC", x"00A9", x"00AD", x"FFA4",
  x"002D", x"0130", x"015F", x"021B"
  );

  signal s_dummy_gyroy_lut : dummy_lut_t := (
  x"0000", x"0000", x"0001", x"0000", x"000D", x"000D", x"0008", x"0024",
  x"0057", x"007B", x"008D", x"0092", x"00EE", x"00EA", x"011B", x"01DC",
  x"0291", x"021C", x"FF5D", x"FD39", x"FD85", x"FE43", x"FEAB", x"FF5F",
  x"FF9A", x"FEA1", x"0FE9", x"FDE6", x"FDDA", x"FE46", x"FE40", x"FE18",
  x"FE5A", x"FE80", x"FE83", x"FDF0", x"FD7F", x"FD68", x"FD98", x"FDC2",
  x"FD16", x"FCED", x"FC50", x"FC62", x"FCDB", x"FD37", x"FCA5", x"FD29",
  x"FDCB", x"FD2B", x"FCE3", x"FDE6", x"FE76", x"FE30", x"FD3F", x"0FD6",
  x"FD47", x"FE64", x"FF51", x"FF4D", x"FE86", x"FE42", x"FE70", x"FE36",
  x"FE74", x"FEF1", x"FF15", x"FE53", x"FD6E", x"FD8C", x"FDDF", x"FEA6",
  x"0FFF", x"FF6B", x"FF54", x"FF76", x"001E", x"00BC", x"01A5", x"022D",
  x"0026", x"0186", x"0095", x"0016", x"00A9", x"001E", x"0088", x"006C",
  x"002E", x"0079", x"012F", x"0319", x"02CA", x"027D", x"017D", x"0215",
  x"0244", x"0277", x"02A3", x"026F", x"0239", x"02C5", x"02B0", x"0277",
  x"0290", x"026B", x"0231", x"0029", x"024C", x"01FF", x"01DA", x"024A",
  x"022A", x"01FB", x"0246", x"0251", x"0212", x"0025", x"0217", x"0214",
  x"023E", x"0221", x"0029", x"01DC", x"01BF", x"0286", x"03B9", x"0324",
  x"0172", x"0069", x"FFA0", x"FF89", x"0033", x"003B", x"008D", x"00B0",
  x"00CA", x"0033", x"FF45", x"FF78", x"FFC2", x"00E6", x"FF5C", x"FC7E",
  x"FC9A", x"FE14", x"FE4E", x"FD74", x"FC35", x"FB39", x"FB4A", x"0FC9",
  x"FCDA", x"FCEE", x"0FD3", x"FDBF", x"FEAE", x"FF5B", x"FFB2", x"FFF6",
  x"FFDE", x"FFC3", x"FFCE", x"004C", x"0094", x"00DD", x"002E", x"029D",
  x"0359", x"03CE", x"0046", x"045F", x"04DC", x"0564", x"0054", x"0447",
  x"043D", x"04CC", x"0535", x"04E1", x"04CB", x"04A8", x"0059", x"05E2",
  x"05AE", x"052E", x"04A1", x"04DA", x"0545", x"0591", x"0632", x"0640",
  x"05CC", x"0610", x"0645", x"0060", x"0679", x"069E", x"0676", x"0068",
  x"05B0", x"05BF", x"0580", x"04B7", x"004A", x"03E7", x"0356", x"02AA",
  x"0274", x"026F", x"0282", x"0295", x"027E", x"01AD", x"00A4", x"FF3F",
  x"FEA3", x"FDF3", x"FCDC", x"0FC8", x"FB19", x"FA60", x"F9C2", x"0FAE",
  x"FA7F", x"F9EE", x"0F97", x"F89A", x"F7AE", x"F6E5", x"F6CD", x"F6D6",
  x"F68F", x"F657", x"F637", x"F670", x"F764", x"F82A", x"F868", x"F8C8",
  x"F8F4", x"F8E2", x"F8FF", x"F936", x"F961", x"F9D5", x"FA8E", x"FACE",
  x"F9EE", x"F8C8", x"F8E5", x"F9A9", x"FA1C", x"FA87", x"FB14", x"FB36",
  x"FAE5", x"FA8A", x"FAE1", x"FB6D", x"FBCA", x"0FC4", x"FC26", x"FC92",
  x"FD22", x"FE33", x"FEE5", x"FEEB", x"FE32", x"FDEB", x"FDF3", x"FDAD",
  x"FCB5", x"FBF1", x"FBD2", x"FC2D", x"FCA6", x"FD24", x"FDB9", x"FEA7",
  x"FF41", x"002E", x"00AB", x"0139", x"0190", x"01E1", x"01F6", x"0251",
  x"034C", x"0430", x"0519", x"05B9", x"05A6", x"054D", x"0551", x"0563",
  x"0544", x"0551", x"05A1", x"0533", x"0462", x"042C", x"0477", x"0477",
  x"0473", x"0429", x"03FA", x"03CF", x"03DB", x"041F", x"04C7", x"04C5",
  x"03F3", x"0337", x"0392", x"03ED", x"038C", x"02CD", x"0029", x"013E",
  x"00F9", x"0017", x"00D2", x"0066", x"003C", x"FFE7", x"FF9A", x"FF38",
  x"0FF7", x"FF13", x"FEFD", x"FEB1", x"FE78", x"FE40", x"FDE4", x"FDEF",
  x"FE4A", x"FEC4", x"FF59", x"FFAD", x"FFF6", x"0076", x"009C", x"007F",
  x"00A2", x"0097", x"0075", x"00AA", x"0113", x"0013", x"00C1", x"0090",
  x"008D", x"0095", x"00D2", x"012C", x"0130", x"00E9", x"00E7", x"00F1",
  x"00FB", x"00ED", x"00B8", x"00C8", x"00CD", x"00B4", x"004E", x"FFDF",
  x"0000", x"0018", x"FFF2", x"FFBF", x"FFBB", x"FF8F", x"FF47", x"0FF2",
  x"FEFE", x"FEF4", x"FEC0", x"FEA2", x"FEA2", x"FE6A", x"FE46", x"FEE8",
  x"FF38", x"FF2B", x"FEDF", x"FED3", x"FEB5", x"FEC7", x"FFA2", x"001B",
  x"FFA3", x"FF2F", x"FEC8", x"FE72", x"FF33", x"0006", x"FFA7", x"FF15",
  x"FF3D", x"003C", x"00B4", x"009E", x"00A4", x"0058", x"0021", x"005D",
  x"00C4", x"001B", x"0156", x"001A", x"0041", x"005F", x"00AC", x"011A",
  x"00FD", x"0070", x"005D", x"00DB", x"0135", x"0015", x"00F2", x"00EC",
  x"00EC", x"0084", x"0014", x"0045", x"00B2", x"0089", x"0014", x"FFFF",
  x"FFEB", x"FFE0", x"FFDD", x"FFED", x"FFF4", x"FFDE", x"FFC9", x"FF8C",
  x"FFB7", x"FFD2", x"FF79", x"FF46", x"FFAD", x"FFFC", x"FFE0", x"FFD3",
  x"FFB8", x"FF83", x"FF4F", x"FF33", x"0FF6", x"FED6", x"FED9", x"FF38",
  x"FF98", x"FFB9", x"FF93", x"FF50", x"FF4A", x"FF82", x"FF9F", x"FFCE",
  x"FFA7", x"FEEC", x"FE1F", x"FD7E", x"FD69", x"FDBF", x"FDA7", x"FCAB",
  x"FBEB", x"FC4B", x"FDDC", x"FEAD", x"FE59", x"FD1E", x"FC4F", x"FC54",
  x"FC3B", x"FC13", x"FBD6", x"FB19", x"FA54", x"FA21", x"FA2A", x"0FA4",
  x"FA1D", x"FA21", x"F9E6", x"FA4F", x"FA44", x"F9CA", x"FAD0", x"FAAA",
  x"FA53", x"FA46", x"FAE2", x"FBDD"
  );

  signal s_dummy_gyroz_lut : dummy_lut_t := (
  x"0001", x"0008", x"000D", x"0009", x"FFFB", x"0FFB", x"000B", x"0040",
  x"003F", x"FFE2", x"0035", x"0051", x"00D4", x"016A", x"015B", x"0135",
  x"023B", x"0266", x"0160", x"00D9", x"FFDF", x"0001", x"0014", x"0038",
  x"0082", x"00B7", x"FF52", x"001E", x"000A", x"0050", x"0049", x"0001",
  x"0025", x"008D", x"0122", x"0145", x"014A", x"014E", x"013C", x"013E",
  x"0131", x"01FC", x"0265", x"0214", x"01EC", x"021D", x"024D", x"023C",
  x"02C8", x"038B", x"0363", x"036E", x"03DF", x"0043", x"046B", x"04AD",
  x"04D5", x"0475", x"03C5", x"0369", x"032D", x"027C", x"0293", x"0319",
  x"037B", x"03C4", x"0382", x"0317", x"02A2", x"0297", x"02ED", x"0428",
  x"049D", x"03F1", x"0350", x"035A", x"0441", x"0539", x"05E6", x"067E",
  x"0660", x"05B1", x"041A", x"0282", x"002E", x"0143", x"016F", x"022B",
  x"0328", x"042E", x"04FD", x"04AC", x"046D", x"0353", x"0295", x"0290",
  x"02C9", x"0293", x"0284", x"0028", x"0195", x"0158", x"0111", x"00A2",
  x"003F", x"FFD3", x"FFA4", x"FF3F", x"FF25", x"FF2C", x"0FF5", x"FEDF",
  x"FE76", x"FE59", x"FE64", x"FE87", x"FEB5", x"FE77", x"FE82", x"FEA4",
  x"FEDE", x"0FFD", x"FF40", x"FF55", x"FF28", x"0FF1", x"000A", x"FF43",
  x"FE87", x"FE9F", x"FEBF", x"FF2C", x"00C5", x"00B1", x"FF35", x"FE90",
  x"FE9D", x"FE99", x"FE75", x"FE8F", x"FF27", x"FF2E", x"FDC7", x"FB6E",
  x"FB7C", x"0FC6", x"FC23", x"FC42", x"FC3C", x"FBB3", x"FB1E", x"FB75",
  x"FBD9", x"FBC0", x"FBA1", x"FC18", x"FC69", x"FCE0", x"FD1C", x"FD66",
  x"FDB7", x"FD80", x"FD2D", x"FD2A", x"FD5C", x"FD97", x"FE1B", x"FECC",
  x"FEC1", x"FE25", x"FDFB", x"0FE7", x"FE5D", x"FEBD", x"FF56", x"FFE3",
  x"00E1", x"01A4", x"018E", x"0168", x"0143", x"0140", x"00E5", x"0055",
  x"0049", x"0088", x"00E9", x"0142", x"0154", x"0175", x"0111", x"0040",
  x"FFBC", x"FFCD", x"000F", x"00A7", x"00FB", x"00E8", x"00A5", x"0037",
  x"0021", x"FFE3", x"FF76", x"FF50", x"FF5A", x"FF2D", x"FEFD", x"FF48",
  x"FFAF", x"FFC0", x"FF84", x"FEC4", x"FE93", x"FEAF", x"FF3B", x"FFE1",
  x"0073", x"00C7", x"00D1", x"00C2", x"0097", x"0078", x"0041", x"004A",
  x"FFFB", x"0040", x"019D", x"0258", x"02C2", x"0213", x"0187", x"011F",
  x"00D3", x"00CB", x"00C6", x"0150", x"01E9", x"0154", x"000E", x"FF70",
  x"FF4A", x"FF4D", x"FF29", x"FEE5", x"FED0", x"FF9D", x"003F", x"FFFA",
  x"FF98", x"FFD0", x"0029", x"00B0", x"00F7", x"00D6", x"0083", x"006B",
  x"00C1", x"015C", x"0116", x"0025", x"FFE6", x"0055", x"00BB", x"00A1",
  x"001F", x"0001", x"FFEC", x"FFF5", x"005E", x"0077", x"0066", x"0056",
  x"008F", x"00EB", x"0014", x"00C9", x"00A5", x"00AE", x"00B5", x"00D4",
  x"0077", x"FFDB", x"FFB8", x"FFC3", x"FFE9", x"FFFC", x"FFB3", x"FF55",
  x"FEFF", x"FEA7", x"FE32", x"FDBC", x"FDA7", x"FE23", x"FE94", x"FE9A",
  x"FE8F", x"FE61", x"FE10", x"FE41", x"FEC4", x"FF10", x"FEDE", x"FECA",
  x"FECE", x"FF25", x"FFB6", x"001D", x"0018", x"0022", x"0048", x"0011",
  x"FFBE", x"FFBF", x"FF9C", x"FF7C", x"FF83", x"FF95", x"FFC9", x"000E",
  x"004E", x"0087", x"0054", x"0002", x"FFFB", x"002C", x"005E", x"0050",
  x"000C", x"FFDD", x"FFE5", x"0015", x"0033", x"0039", x"FFD0", x"FFD5",
  x"FFF5", x"000A", x"0097", x"00A8", x"0064", x"004C", x"003C", x"0069",
  x"0095", x"0043", x"000F", x"0052", x"0097", x"0076", x"0055", x"0041",
  x"0043", x"0027", x"006E", x"007A", x"004C", x"0057", x"00A1", x"00AC",
  x"004A", x"FFAD", x"FFA4", x"FFDA", x"0022", x"005A", x"0049", x"009B",
  x"00B4", x"0068", x"005D", x"00AC", x"0091", x"0048", x"004D", x"0011",
  x"FFFE", x"FFC7", x"FFBF", x"FFA2", x"FF71", x"FF1E", x"FEBA", x"FEBD",
  x"FF15", x"FF44", x"FF17", x"FF3B", x"FF29", x"FECD", x"FE7B", x"FEBF",
  x"FF89", x"FF9C", x"FF55", x"FED4", x"FF11", x"FF70", x"FF3F", x"FEEF",
  x"FF61", x"000D", x"005C", x"003A", x"FFEE", x"FF77", x"FF87", x"FFC0",
  x"FF8E", x"FF40", x"FEBD", x"FEA3", x"FE64", x"FEE7", x"FF81", x"FFEA",
  x"FFC0", x"FF94", x"FFA2", x"0029", x"006B", x"0023", x"0026", x"008F",
  x"0121", x"0188", x"015C", x"0117", x"0183", x"021D", x"022F", x"022A",
  x"01F5", x"01E6", x"01ED", x"021C", x"0246", x"01D4", x"01A9", x"015F",
  x"00E8", x"00D4", x"00E1", x"0090", x"0000", x"0003", x"FFEE", x"FFD0",
  x"FF77", x"0FFC", x"FEDD", x"FEC9", x"FEAA", x"FEA3", x"FE5C", x"FE37",
  x"FE24", x"FD93", x"0FDA", x"FCBB", x"FCEA", x"FD3C", x"FD64", x"FDE2",
  x"FE89", x"FF1C", x"FF89", x"0030", x"00C0", x"011B", x"019C", x"029B",
  x"003E", x"0297", x"0174", x"00A6", x"008B", x"00DB", x"012A", x"013B",
  x"0138", x"00F7", x"00ED", x"011B", x"0087", x"FFF6", x"FFA8", x"FFD5",
  x"0006", x"FFD7", x"FF85", x"FF5A", x"FF45", x"FED1", x"FE98", x"FF2B",
  x"FF7E", x"FF93", x"FF23", x"FF1C"
  );

  signal s_dummy_magx_lut : dummy_lut_t := (
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000"
  );

  signal s_dummy_magy_lut : dummy_lut_t := (
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000"
  );

  signal s_dummy_magz_lut : dummy_lut_t := (
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
  x"0000", x"0000", x"0000", x"0000"
  );

  signal s_dummy_temp_lut : dummy_lut_t := (
  x"0DA0", x"0DA0", x"0DD0", x"0DA0", x"0D70", x"0DA0", x"0DD0", x"0DC0",
  x"0D90", x"0D90", x"0D60", x"00E0", x"0D50", x"0DD0", x"0D90", x"0DA0",
  x"0DC0", x"0DA0", x"0D70", x"0DA0", x"0DE0", x"0DE0", x"00E0", x"0D70",
  x"0DD0", x"0D50", x"0D70", x"00E0", x"0DC0", x"0DA0", x"0DA0", x"0DE0",
  x"0D60", x"0DA0", x"0D90", x"0DA0", x"0DC0", x"00E0", x"0D60", x"0DE0",
  x"0D70", x"0D70", x"0DA0", x"0DC0", x"0E10", x"0DA0", x"0D90", x"0DD0",
  x"0DC0", x"0DD0", x"0DD0", x"0DA0", x"0D70", x"0DA0", x"0D90", x"0DE0",
  x"00E0", x"0DD0", x"0DA0", x"0D50", x"0DC0", x"0DE0", x"0DA0", x"0DA0",
  x"0D30", x"0E10", x"00E0", x"0D60", x"00E0", x"0DA0", x"0D90", x"0DA0",
  x"0DA0", x"0DA0", x"0D70", x"0DC0", x"00E0", x"0D50", x"0DD0", x"0DA0",
  x"0DA0", x"0DC0", x"0DD0", x"0D90", x"0DA0", x"0D50", x"0DD0", x"0E10",
  x"0D90", x"0DD0", x"0D70", x"0DA0", x"0DC0", x"0DA0", x"0DA0", x"0DC0",
  x"0DC0", x"0DC0", x"0D70", x"00E0", x"00E0", x"0DA0", x"0D70", x"0D60",
  x"0DC0", x"0DC0", x"0D60", x"0DD0", x"0D60", x"0DA0", x"0D50", x"0D50",
  x"0DD0", x"00E0", x"0DD0", x"0DE0", x"0DA0", x"0DD0", x"0DC0", x"0D90",
  x"0DE0", x"0DA0", x"0DC0", x"0DC0", x"0D70", x"0DE0", x"0DE0", x"0DA0",
  x"0DE0", x"0DA0", x"0D60", x"0DA0", x"0DC0", x"0DD0", x"0DC0", x"0D90",
  x"0DE0", x"0DA0", x"0E10", x"0D90", x"0DA0", x"0DA0", x"0D70", x"0DA0",
  x"0E10", x"0DC0", x"0DA0", x"0DA0", x"00E0", x"0D90", x"0DA0", x"0DC0",
  x"0DE0", x"0DA0", x"0DC0", x"0D50", x"0DA0", x"00E0", x"0DA0", x"0DC0",
  x"00E0", x"0DE0", x"0DA0", x"0D90", x"0DD0", x"0DA0", x"0DA0", x"0DA0",
  x"0D70", x"0DD0", x"0D70", x"0DA0", x"00E0", x"0D90", x"0DC0", x"0DA0",
  x"0D50", x"0DA0", x"00E0", x"0DA0", x"0DA0", x"0DE0", x"0DA0", x"0DA0",
  x"0D60", x"0DA0", x"0DA0", x"0DA0", x"0DC0", x"0DA0", x"0DA0", x"0DA0",
  x"0DD0", x"0DA0", x"0DA0", x"0DA0", x"0DE0", x"0DA0", x"0DD0", x"0DC0",
  x"0DC0", x"0DC0", x"0D70", x"0DC0", x"0DD0", x"0D60", x"0DA0", x"0D70",
  x"0D60", x"0DA0", x"0DC0", x"0DA0", x"0DC0", x"0D70", x"0DA0", x"0D30",
  x"0DA0", x"0DA0", x"0DA0", x"0DC0", x"0D90", x"0DC0", x"0DC0", x"0D90",
  x"0DA0", x"0D50", x"0DE0", x"0DC0", x"0DC0", x"0DD0", x"0DA0", x"0DA0",
  x"0D70", x"0D50", x"0DC0", x"0DD0", x"0DA0", x"0DD0", x"0D50", x"0DE0",
  x"0DC0", x"0DD0", x"0DA0", x"0DC0", x"0DA0", x"0DE0", x"0D50", x"00E0",
  x"0D90", x"0DD0", x"0D70", x"0D70", x"0DA0", x"0DA0", x"0E10", x"0DE0",
  x"0DD0", x"0DA0", x"0D60", x"0D70", x"0DC0", x"0DA0", x"0DA0", x"0D70",
  x"0D60", x"0DA0", x"0DD0", x"0DD0", x"0D90", x"0DA0", x"0DA0", x"00E0",
  x"0DD0", x"0E10", x"0D90", x"0DD0", x"0D90", x"0D70", x"0DA0", x"0DE0",
  x"0DE0", x"0D50", x"0DA0", x"0DA0", x"0DA0", x"0D50", x"0DC0", x"0DD0",
  x"0D60", x"0DA0", x"0D90", x"0DA0", x"0DD0", x"0E10", x"0DD0", x"0D90",
  x"0DD0", x"0DA0", x"0D70", x"0DE0", x"0DA0", x"0D70", x"0DC0", x"0DC0",
  x"00E0", x"0DC0", x"0DD0", x"0DA0", x"0DE0", x"0DE0", x"00E0", x"0DA0",
  x"00E0", x"0DA0", x"0DA0", x"0D70", x"0DA0", x"0D70", x"0DA0", x"0DC0",
  x"0DD0", x"0D70", x"0D90", x"0DC0", x"0D60", x"0DC0", x"0DD0", x"00E0",
  x"0DC0", x"0D60", x"0DC0", x"0DA0", x"0DA0", x"0DA0", x"0D30", x"0DE0",
  x"0D70", x"0DE0", x"0DE0", x"0D60", x"0DA0", x"0DC0", x"0D50", x"0DA0",
  x"0DD0", x"0D70", x"0D60", x"0D70", x"0D90", x"0DC0", x"0DA0", x"00E0",
  x"0D60", x"0DC0", x"0DC0", x"0DE0", x"0DD0", x"0D50", x"0DE0", x"0DA0",
  x"0D90", x"0DD0", x"0DD0", x"0D70", x"0DD0", x"0D70", x"0DC0", x"0DA0",
  x"0DC0", x"0DA0", x"0D70", x"0DA0", x"0E10", x"0E10", x"0DC0", x"0D90",
  x"0D70", x"0DE0", x"0DA0", x"0DC0", x"0DA0", x"00E0", x"0DA0", x"0D70",
  x"0DA0", x"0DC0", x"00E0", x"0D70", x"0D70", x"00E0", x"0DA0", x"0DD0",
  x"0DE0", x"0D70", x"0DD0", x"0DD0", x"0D70", x"0DD0", x"0DC0", x"00E0",
  x"0DD0", x"0D70", x"0DC0", x"0DE0", x"0DC0", x"0D70", x"0D90", x"0DD0",
  x"0D90", x"0D70", x"0DA0", x"0DC0", x"0DA0", x"0DE0", x"0D90", x"0DC0",
  x"0DD0", x"0DE0", x"0DC0", x"0D60", x"00E0", x"0E10", x"0D60", x"0DD0",
  x"0DA0", x"0DE0", x"0DE0", x"0D60", x"00E0", x"0DE0", x"0D90", x"0DD0",
  x"0D70", x"0DA0", x"00E0", x"0D70", x"0DA0", x"0DC0", x"0DC0", x"0DC0",
  x"0D70", x"0DC0", x"0DD0", x"0D70", x"0DE0", x"0D70", x"0D70", x"0DD0",
  x"0D50", x"0DD0", x"0DE0", x"00E0", x"0DC0", x"0D60", x"0DC0", x"0DA0",
  x"0DA0", x"0DC0", x"0D70", x"0DD0", x"0D60", x"0DD0", x"0DC0", x"0DC0",
  x"0DD0", x"0DC0", x"0D70", x"0DC0", x"0DC0", x"0DC0", x"00E0", x"0DD0",
  x"0DD0", x"00E0", x"0DA0", x"0DA0", x"0DC0", x"0D90", x"0DD0", x"0D90",
  x"0DD0", x"0D60", x"0DA0", x"0D90", x"0DA0", x"0DC0", x"0DA0", x"0DC0",
  x"0DC0", x"0DA0", x"0DE0", x"0DA0", x"0D90", x"0DA0", x"0DA0", x"0DD0",
  x"00E0", x"0D30", x"00E0", x"0D90"
  );
  -- Counter to keep track of the current index in the LUT
  signal s_index_cnt : integer range 0 to G_IMU_DATA_CNT - 1 := 0;

begin

  -- Process to increment the index used for the luts
  P_switching_luts : process (clk_i, rst_i)
  begin
    if rst_i = '1' then
      s_index_cnt <= 0;
    elsif clk_i'event and clk_i = '1' then
      if tick_i = '1' then
        if s_index_cnt < G_IMU_DATA_CNT - 1 then
          s_index_cnt <= s_index_cnt + 1;
        else
          s_index_cnt <= 0;
        end if;
      end if;
    end if;
  end process;

  -- Output the value from the lookup table based on the index
  accel_xout_o <= s_dummy_accelx_lut(s_index_cnt);
  accel_yout_o <= s_dummy_accely_lut(s_index_cnt);
  accel_zout_o <= s_dummy_accelz_lut(s_index_cnt);
  gyro_xout_o  <= s_dummy_gyrox_lut(s_index_cnt);
  gyro_yout_o  <= s_dummy_gyroy_lut(s_index_cnt);
  gyro_zout_o  <= s_dummy_gyroz_lut(s_index_cnt);
  mag_xout_o   <= s_dummy_magx_lut(s_index_cnt);
  mag_yout_o   <= s_dummy_magy_lut(s_index_cnt);
  mag_zout_o   <= s_dummy_magz_lut(s_index_cnt);
  temp_out_o   <= s_dummy_temp_lut(s_index_cnt);
end architecture;
